module Somador4b(
    input logic[3:0] a, b,
    output logic[3:0] s);

    assign s = a + b;

endmodule
